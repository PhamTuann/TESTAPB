`ifndef PAC
`define PAC

class Packet;
	rand reg [7:0] PWDATA;
endclass

`endif 